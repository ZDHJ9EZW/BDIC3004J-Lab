module A(output [7:0] ALU_out, input [7:0] Data_A, Data_B, input [2:0] Opcode);
	
	Lab1 M1 (ALU_out, Data_A, Data_B, Opcode);
endmodule